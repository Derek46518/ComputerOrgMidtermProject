`timescale 1ns/1ns
module Multiplier( clk, dataA, dataB, Signal, dataOut, reset);
input clk, reset;
input [31:0] dataA, dataB;
input [5:0] Signal;
output[63:0] dataOut;
reg[63:0] Product,temp;
reg[31:0] B;
parameter MULTU=6'b011001;
parameter OUT = 6'b111111;

always@(posedge clk or reset)
    begin
        if (reset) 
        begin
            assign Product = 64'b0;
            assign temp = {32'b0,dataA[31:0]};
            assign B={dataB[31:0]};
        end
    
        else
        begin
        case ( Signal )
  		MULTU:
		begin
            if(B[0]) begin
                assign Product = temp+Product;
            end

            assign B = B >> 1;
            assign temp = temp << 1;
		end
  		OUT:
		begin
			Product <= 64'b0;
            temp <= {32'b0,dataA[31:0]};
            B <={dataB[31:0]};
        end
		
		endcase
        end
        
    end
assign dataOut = Product;
endmodule